package in_out_matrix is
    
    TYPE in_array is ARRAY  (natural range <>) of std_logic_vector(7 downto 0);
    TYPE tf_array is ARRAY  (natural range <>) of std_logic_vector(7 downto 0);  
    TYPE out_array is ARRAY (natural range <>) of std_logic_vector(7 downto 0); 

end package; 