-------------------------------------------
-- Project			: ELEC562 32 BIT FFT 
-- Author			: Matthew Stein
-- Date				: 2019-04-22
-- File				: single_dft_tb.vhd
-- Description		: Test bench for stage2. 
--                    Twiddle factors are assuemd to be accurate and included as inputs. 
-- 
-------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use work.in_out_matrix.all;

entity single_dft_tb is
end single_dft_tb;

architecture test of single_dft_tb is 
  
    signal real_in_s                : in_array(0 to 1); 
    signal imag_in_s                : in_array(0 to 1); 
    signal tf_real_s                : std_logic_vector(15 downto 0);
    signal tf_imag_s                : std_logic_vector(15 downto 0);
    signal real_out_s               : out_array(0 to 1); 
    signal imag_out_s               : out_array(0 to 1); 
    signal rst_s                    : std_logic; 
    -- Clocks 
    signal clk_s                    : std_logic; 
    constant clock_period           : time := 10 ns; 

    begin
        single_dft_tb : entity work.single_dft(structural)
        port map(
            real_in => real_in_s, 
            imag_in => imag_in_s, 
            tf_real => tf_real_s, 
            tf_imag => tf_imag_s, 
            real_out => real_out_s, 
            imag_out => imag_out_s, 
            rst => rst_s, 
            clk => clk_s
        );

    clock_process : process
    begin
        clk_s <= '0';
        wait for clock_period/2;
        clk_s <= '1';
        wait for clock_period/2;
    end process;
    
    -- Note: One clock cycle is set to 10s, and each Single DFT block takes 2 clock cycles.
    -- Recall: Inputs must be constrained to a value only using 11 bits of the input (for growth) 
            -- Thus Inputs must be less than or equal to x"07ff" 
    stim_proc : process
        begin
            wait for 20 ns;
            rst_s <= '1'; 
            wait for 20 ns; 
            rst_s <= '0'; 
            wait for 20 ns; 

          
            tf_real_s <=  ( x"7fff");
            tf_imag_s <=  ( x"0000");
        
            real_in_s <= (x"0000",x"0001");
            imag_in_s <= (x"0000",x"0001");

            wait for 20 ns;
            
            real_in_s <= (x"0001",x"0000");

            imag_in_s <= (x"0001",x"0000");
            
            wait for 20 ns;
            rst_s <= '1'; 
            wait for 20 ns; 
            rst_s <= '0';
            
            tf_real_s <=  ( x"7D8A");
            tf_imag_s <=  ( x"18F9");
            
            real_in_s <= (x"0000",x"0001");
            imag_in_s <= (x"0000",x"0001");
           
            wait for 20 ns;
                       
            real_in_s <= (x"0001",x"0000");          
            imag_in_s <= (x"0001",x"0000");
            
            wait for 20 ns; 
            rst_s <= '0'; 
            wait for 20 ns; 
            

        end process;


    end test;


